** Generated for: hspiceD
** Generated on: Dec  7 12:58:19 2024
** Design library name: trail
** Design cell name: AND
** Design view name: schematic



** Library name: trail
** Cell name: AND
** View name: schematic
xm4 y net1 gnd gnd nch_lvt_mac l=16e-9 nfin=1 w=10e-9 multi=1 nf=1 sa=90e-9 sb=90e-9
xm1 net2 b gnd gnd nch_lvt_mac l=16e-9 nfin=2 w=58e-9 multi=1 nf=1 sa=90e-9 sb=90e-9
xm0 net1 a net2 gnd nch_lvt_mac l=16e-9 nfin=2 w=58e-9 multi=1 nf=1 sa=90e-9 sb=90e-9
xm5 y net1 vdd vdd pch_lvt_mac l=16e-9 nfin=1 w=10e-9 multi=1 nf=1 sa=90e-9 sb=90e-9
xm3 net1 b vdd vdd pch_lvt_mac l=16e-9 nfin=1 w=10e-9 multi=1 nf=1 sa=90e-9 sb=90e-9
xm2 net1 a vdd vdd pch_lvt_mac l=16e-9 nfin=1 w=10e-9 multi=1 nf=1 sa=90e-9 sb=90e-9
.END

